module picmicro_midrange_core_de2_115(
	input wire CLOCK_50
);

//this implementation will mimic the 16f628a


endmodule

