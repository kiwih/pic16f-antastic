module instruction_decoder(
	input wire clk,
	
	input wire [13:0] instr_current,
	
	output wire instr_rd_en
);



endmodule
