module picmicro_midrange_core_de2_115(
	input wire CLOCK_50
);


endmodule

