localparam portb_address	=		9'bz00000110;
localparam trisb_address	=		9'bz10000110;

localparam porta_address	=		9'h05;
localparam trisa_address	=		9'h85;

localparam txsta_address 	=		9'h98;
localparam spbrg_address	=		9'h99;
localparam rcsta_address	=		9'h18;
localparam txreg_address	=		9'h19;
localparam rcreg_address	=		9'h1a;