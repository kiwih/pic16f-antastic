module picmicro_midrange_core(
	input wire clk
);

endmodule
