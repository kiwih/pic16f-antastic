localparam portb_address	=		9'bz00000110;
localparam trisb_address	=		9'bz10000110;

localparam porta_address	=		9'h05;
localparam trisa_address	=		9'h85;



